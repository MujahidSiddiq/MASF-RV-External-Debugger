`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/23/2024 12:06:19 PM
// Design Name: 
// Module Name: mux_2x1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux_2x1(

    input  logic              select,
    input  logic [31:0]       data0,
    input  logic [31:0]       data1,
    output logic [31:0]       out
    
    
    );
    
    assign out = select ? data1 :  data0;

    
endmodule
