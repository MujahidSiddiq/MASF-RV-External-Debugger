`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/23/2024 12:09:24 PM
// Design Name: 
// Module Name: Plus_4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Plus_4(

     input  logic [31:0]     in,
     output logic [31:0]     out

    );

    assign out     =         in + 4 ;

    
endmodule
